// Code your design here
`include "programCounter.v"
`include "mux2to1.v"
`include "instructionMemory.v"
`include "instructionParser.v"
`include "dataGenerator.v"
`include "adder.v"
`include "ALU_64_bit.v"
`include "ALUcontrol.v"
`include "controlUnit.v"
`include "dataMemory.v"
`include "registerFile.v"
`include "singleProcessor.v"